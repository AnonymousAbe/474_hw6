module tas(
	


);



endmodule
